library verilog;
use verilog.vl_types.all;
entity lcd_driver_vlg_vec_tst is
end lcd_driver_vlg_vec_tst;
