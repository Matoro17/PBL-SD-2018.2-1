library verilog;
use verilog.vl_types.all;
entity Nios_mm_interconnect_0 is
    port(
        Clk_clk_clk     : in     vl_logic;
        Nios_reset_n_reset_bridge_in_reset_reset: in     vl_logic;
        Nios_data_master_address: in     vl_logic_vector(15 downto 0);
        Nios_data_master_waitrequest: out    vl_logic;
        Nios_data_master_byteenable: in     vl_logic_vector(3 downto 0);
        Nios_data_master_read: in     vl_logic;
        Nios_data_master_readdata: out    vl_logic_vector(31 downto 0);
        Nios_data_master_write: in     vl_logic;
        Nios_data_master_writedata: in     vl_logic_vector(31 downto 0);
        Nios_data_master_debugaccess: in     vl_logic;
        Nios_instruction_master_address: in     vl_logic_vector(15 downto 0);
        Nios_instruction_master_waitrequest: out    vl_logic;
        Nios_instruction_master_read: in     vl_logic;
        Nios_instruction_master_readdata: out    vl_logic_vector(31 downto 0);
        dip_0_s1_address: out    vl_logic_vector(1 downto 0);
        dip_0_s1_readdata: in     vl_logic_vector(31 downto 0);
        dip_1_s1_address: out    vl_logic_vector(1 downto 0);
        dip_1_s1_readdata: in     vl_logic_vector(31 downto 0);
        dip_2_s1_address: out    vl_logic_vector(1 downto 0);
        dip_2_s1_readdata: in     vl_logic_vector(31 downto 0);
        dip_3_s1_address: out    vl_logic_vector(1 downto 0);
        dip_3_s1_readdata: in     vl_logic_vector(31 downto 0);
        Jtag_avalon_jtag_slave_address: out    vl_logic_vector(0 downto 0);
        Jtag_avalon_jtag_slave_write: out    vl_logic;
        Jtag_avalon_jtag_slave_read: out    vl_logic;
        Jtag_avalon_jtag_slave_readdata: in     vl_logic_vector(31 downto 0);
        Jtag_avalon_jtag_slave_writedata: out    vl_logic_vector(31 downto 0);
        Jtag_avalon_jtag_slave_waitrequest: in     vl_logic;
        Jtag_avalon_jtag_slave_chipselect: out    vl_logic;
        led_1_s1_address: out    vl_logic_vector(1 downto 0);
        led_1_s1_write  : out    vl_logic;
        led_1_s1_readdata: in     vl_logic_vector(31 downto 0);
        led_1_s1_writedata: out    vl_logic_vector(31 downto 0);
        led_1_s1_chipselect: out    vl_logic;
        led_2_s1_address: out    vl_logic_vector(1 downto 0);
        led_2_s1_write  : out    vl_logic;
        led_2_s1_readdata: in     vl_logic_vector(31 downto 0);
        led_2_s1_writedata: out    vl_logic_vector(31 downto 0);
        led_2_s1_chipselect: out    vl_logic;
        led_3_s1_address: out    vl_logic_vector(1 downto 0);
        led_3_s1_write  : out    vl_logic;
        led_3_s1_readdata: in     vl_logic_vector(31 downto 0);
        led_3_s1_writedata: out    vl_logic_vector(31 downto 0);
        led_3_s1_chipselect: out    vl_logic;
        led_4_s1_address: out    vl_logic_vector(1 downto 0);
        led_4_s1_write  : out    vl_logic;
        led_4_s1_readdata: in     vl_logic_vector(31 downto 0);
        led_4_s1_writedata: out    vl_logic_vector(31 downto 0);
        led_4_s1_chipselect: out    vl_logic;
        led_5_s1_address: out    vl_logic_vector(1 downto 0);
        led_5_s1_write  : out    vl_logic;
        led_5_s1_readdata: in     vl_logic_vector(31 downto 0);
        led_5_s1_writedata: out    vl_logic_vector(31 downto 0);
        led_5_s1_chipselect: out    vl_logic;
        memory_s1_address: out    vl_logic_vector(11 downto 0);
        memory_s1_write : out    vl_logic;
        memory_s1_readdata: in     vl_logic_vector(31 downto 0);
        memory_s1_writedata: out    vl_logic_vector(31 downto 0);
        memory_s1_byteenable: out    vl_logic_vector(3 downto 0);
        memory_s1_chipselect: out    vl_logic;
        memory_s1_clken : out    vl_logic;
        Nios_jtag_debug_module_address: out    vl_logic_vector(8 downto 0);
        Nios_jtag_debug_module_write: out    vl_logic;
        Nios_jtag_debug_module_read: out    vl_logic;
        Nios_jtag_debug_module_readdata: in     vl_logic_vector(31 downto 0);
        Nios_jtag_debug_module_writedata: out    vl_logic_vector(31 downto 0);
        Nios_jtag_debug_module_byteenable: out    vl_logic_vector(3 downto 0);
        Nios_jtag_debug_module_waitrequest: in     vl_logic;
        Nios_jtag_debug_module_debugaccess: out    vl_logic;
        pushbutton_1_s1_address: out    vl_logic_vector(1 downto 0);
        pushbutton_1_s1_write: out    vl_logic;
        pushbutton_1_s1_readdata: in     vl_logic_vector(31 downto 0);
        pushbutton_1_s1_writedata: out    vl_logic_vector(31 downto 0);
        pushbutton_1_s1_chipselect: out    vl_logic;
        pushbutton_2_s1_address: out    vl_logic_vector(1 downto 0);
        pushbutton_2_s1_write: out    vl_logic;
        pushbutton_2_s1_readdata: in     vl_logic_vector(31 downto 0);
        pushbutton_2_s1_writedata: out    vl_logic_vector(31 downto 0);
        pushbutton_2_s1_chipselect: out    vl_logic
    );
end Nios_mm_interconnect_0;
