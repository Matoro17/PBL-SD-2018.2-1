library verilog;
use verilog.vl_types.all;
entity Nios_Nios_nios2_performance_monitors is
end Nios_Nios_nios2_performance_monitors;
